module adder (input [1:0] a, input [1:0] b, output [1:0] y);
    assign y = a + b;
endmodule